// Video_System.v


`timescale 1 ps / 1 ps
module Video_System (
		output wire        VGA_CLK_from_the_VGA_Controller,                     //   VGA_Controller_external_interface.CLK
		output wire        VGA_HS_from_the_VGA_Controller,                      //                                    .HS
		output wire        VGA_VS_from_the_VGA_Controller,                      //                                    .VS
		output wire        VGA_BLANK_from_the_VGA_Controller,                   //                                    .BLANK
		output wire        VGA_SYNC_from_the_VGA_Controller,                    //                                    .SYNC
		output wire [7:0]  VGA_R_from_the_VGA_Controller,                       //                                    .R
		output wire [7:0]  VGA_G_from_the_VGA_Controller,                       //                                    .G
		output wire [7:0]  VGA_B_from_the_VGA_Controller,                       //                                    .B
		input  wire        reset_n,                                             //                    clk_clk_in_reset.reset_n
		inout  wire        I2C_SDAT_to_and_from_the_AV_Config,                  //        AV_Config_external_interface.SDAT
		output wire        I2C_SCLK_from_the_AV_Config,                         //                                    .SCLK
		input  wire        clk,                                                 //                          clk_clk_in.clk
		inout  wire [15:0] SRAM_DQ_to_and_from_the_Pixel_Buffer,                //     Pixel_Buffer_external_interface.DQ
		output wire [19:0] SRAM_ADDR_from_the_Pixel_Buffer,                     //                                    .ADDR
		output wire        SRAM_LB_N_from_the_Pixel_Buffer,                     //                                    .LB_N
		output wire        SRAM_UB_N_from_the_Pixel_Buffer,                     //                                    .UB_N
		output wire        SRAM_CE_N_from_the_Pixel_Buffer,                     //                                    .CE_N
		output wire        SRAM_OE_N_from_the_Pixel_Buffer,                     //                                    .OE_N
		output wire        SRAM_WE_N_from_the_Pixel_Buffer,                     //                                    .WE_N
		input  wire        Video_In_Decoder_external_interface_PIXEL_CLK,       // Video_In_Decoder_external_interface.PIXEL_CLK
		input  wire        Video_In_Decoder_external_interface_LINE_VALID,      //                                    .LINE_VALID
		input  wire        Video_In_Decoder_external_interface_FRAME_VALID,     //                                    .FRAME_VALID
		input  wire        Video_In_Decoder_external_interface_pixel_clk_reset, //                                    .pixel_clk_reset
		input  wire [9:0]  Video_In_Decoder_external_interface_PIXEL_DATA       //                                    .PIXEL_DATA
	);

	wire         pixel_scaler_avalon_scaler_source_endofpacket;                                                              // Pixel_Scaler:stream_out_endofpacket -> Dual_Clock_FIFO:stream_in_endofpacket
	wire         pixel_scaler_avalon_scaler_source_valid;                                                                    // Pixel_Scaler:stream_out_valid -> Dual_Clock_FIFO:stream_in_valid
	wire         pixel_scaler_avalon_scaler_source_startofpacket;                                                            // Pixel_Scaler:stream_out_startofpacket -> Dual_Clock_FIFO:stream_in_startofpacket
	wire  [29:0] pixel_scaler_avalon_scaler_source_data;                                                                     // Pixel_Scaler:stream_out_data -> Dual_Clock_FIFO:stream_in_data
	wire         pixel_scaler_avalon_scaler_source_ready;                                                                    // Dual_Clock_FIFO:stream_in_ready -> Pixel_Scaler:stream_out_ready
	wire         pixel_rgb_resampler_avalon_rgb_source_endofpacket;                                                          // Pixel_RGB_Resampler:stream_out_endofpacket -> Pixel_Scaler:stream_in_endofpacket
	wire         pixel_rgb_resampler_avalon_rgb_source_valid;                                                                // Pixel_RGB_Resampler:stream_out_valid -> Pixel_Scaler:stream_in_valid
	wire         pixel_rgb_resampler_avalon_rgb_source_startofpacket;                                                        // Pixel_RGB_Resampler:stream_out_startofpacket -> Pixel_Scaler:stream_in_startofpacket
	wire  [29:0] pixel_rgb_resampler_avalon_rgb_source_data;                                                                 // Pixel_RGB_Resampler:stream_out_data -> Pixel_Scaler:stream_in_data
	wire         pixel_rgb_resampler_avalon_rgb_source_ready;                                                                // Pixel_Scaler:stream_in_ready -> Pixel_RGB_Resampler:stream_out_ready
	wire         pixel_buffer_dma_avalon_pixel_source_endofpacket;                                                           // Pixel_Buffer_DMA:stream_endofpacket -> Pixel_RGB_Resampler:stream_in_endofpacket
	wire         pixel_buffer_dma_avalon_pixel_source_valid;                                                                 // Pixel_Buffer_DMA:stream_valid -> Pixel_RGB_Resampler:stream_in_valid
	wire         pixel_buffer_dma_avalon_pixel_source_startofpacket;                                                         // Pixel_Buffer_DMA:stream_startofpacket -> Pixel_RGB_Resampler:stream_in_startofpacket
	wire  [15:0] pixel_buffer_dma_avalon_pixel_source_data;                                                                  // Pixel_Buffer_DMA:stream_data -> Pixel_RGB_Resampler:stream_in_data
	wire         pixel_buffer_dma_avalon_pixel_source_ready;                                                                 // Pixel_RGB_Resampler:stream_in_ready -> Pixel_Buffer_DMA:stream_ready
	wire         dual_clock_fifo_avalon_dc_buffer_source_endofpacket;                                                        // Dual_Clock_FIFO:stream_out_endofpacket -> VGA_Controller:endofpacket
	wire         dual_clock_fifo_avalon_dc_buffer_source_valid;                                                              // Dual_Clock_FIFO:stream_out_valid -> VGA_Controller:valid
	wire         dual_clock_fifo_avalon_dc_buffer_source_startofpacket;                                                      // Dual_Clock_FIFO:stream_out_startofpacket -> VGA_Controller:startofpacket
	wire  [29:0] dual_clock_fifo_avalon_dc_buffer_source_data;                                                               // Dual_Clock_FIFO:stream_out_data -> VGA_Controller:data
	wire         dual_clock_fifo_avalon_dc_buffer_source_ready;                                                              // VGA_Controller:ready -> Dual_Clock_FIFO:stream_out_ready
	wire         video_rgb_resampler_avalon_rgb_source_endofpacket;                                                          // Video_RGB_Resampler:stream_out_endofpacket -> Video_Clipper:stream_in_endofpacket
	wire         video_rgb_resampler_avalon_rgb_source_valid;                                                                // Video_RGB_Resampler:stream_out_valid -> Video_Clipper:stream_in_valid
	wire         video_rgb_resampler_avalon_rgb_source_startofpacket;                                                        // Video_RGB_Resampler:stream_out_startofpacket -> Video_Clipper:stream_in_startofpacket
	wire  [15:0] video_rgb_resampler_avalon_rgb_source_data;                                                                 // Video_RGB_Resampler:stream_out_data -> Video_Clipper:stream_in_data
	wire         video_rgb_resampler_avalon_rgb_source_ready;                                                                // Video_Clipper:stream_in_ready -> Video_RGB_Resampler:stream_out_ready
	wire         video_clipper_avalon_clipper_source_endofpacket;                                                            // Video_Clipper:stream_out_endofpacket -> Video_Scaler:stream_in_endofpacket
	wire         video_clipper_avalon_clipper_source_valid;                                                                  // Video_Clipper:stream_out_valid -> Video_Scaler:stream_in_valid
	wire         video_clipper_avalon_clipper_source_startofpacket;                                                          // Video_Clipper:stream_out_startofpacket -> Video_Scaler:stream_in_startofpacket
	wire  [15:0] video_clipper_avalon_clipper_source_data;                                                                   // Video_Clipper:stream_out_data -> Video_Scaler:stream_in_data
	wire         video_clipper_avalon_clipper_source_ready;                                                                  // Video_Scaler:stream_in_ready -> Video_Clipper:stream_out_ready
	wire         video_scaler_avalon_scaler_source_endofpacket;                                                              // Video_Scaler:stream_out_endofpacket -> Video_DMA:stream_endofpacket
	wire         video_scaler_avalon_scaler_source_valid;                                                                    // Video_Scaler:stream_out_valid -> Video_DMA:stream_valid
	wire         video_scaler_avalon_scaler_source_startofpacket;                                                            // Video_Scaler:stream_out_startofpacket -> Video_DMA:stream_startofpacket
	wire  [15:0] video_scaler_avalon_scaler_source_data;                                                                     // Video_Scaler:stream_out_data -> Video_DMA:stream_data
	wire         video_scaler_avalon_scaler_source_ready;                                                                    // Video_DMA:stream_ready -> Video_Scaler:stream_out_ready
	wire         clock_signals_sys_clk_clk;                                                                                  // Clock_Signals:sys_clk -> [AV_Config:clk, AV_Config_avalon_av_config_slave_translator:clk, AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:clk, AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, CPU:clk, CPU_data_master_translator:clk, CPU_data_master_translator_avalon_universal_master_0_agent:clk, CPU_instruction_master_translator:clk, CPU_instruction_master_translator_avalon_universal_master_0_agent:clk, CPU_jtag_debug_module_translator:clk, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Dual_Clock_FIFO:clk_stream_in, Onchip_Memory:clk, Onchip_Memory_s1_translator:clk, Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:clk, Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Pixel_Buffer:clk, Pixel_Buffer_DMA:clk, Pixel_Buffer_DMA_avalon_control_slave_translator:clk, Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:clk, Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:clk, Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:clk, Pixel_Buffer_avalon_sram_slave_translator:clk, Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:clk, Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Pixel_RGB_Resampler:clk, Pixel_Scaler:clk, Video_Clipper:clk, Video_DMA:clk, Video_DMA_avalon_dma_control_slave_translator:clk, Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:clk, Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Video_DMA_avalon_dma_master_translator:clk, Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:clk, Video_In_Decoder:clk, Video_RGB_Resampler:clk, Video_Scaler:clk, addr_router:clk, addr_router_001:clk, addr_router_002:clk, addr_router_003:clk, burst_adapter:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_demux_003:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, irq_mapper:clk, limiter:clk, limiter_001:clk, limiter_002:clk, limiter_003:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, width_adapter:clk, width_adapter_001:clk]
	wire         clock_signals_vga_clk_clk;                                                                                  // Clock_Signals:VGA_CLK -> [Dual_Clock_FIFO:clk_stream_out, VGA_Controller:clk, rst_controller_001:clk]
	wire         video_in_decoder_avalon_decoder_source_endofpacket;                                                         // Video_In_Decoder:stream_out_endofpacket -> Video_RGB_Resampler:stream_in_endofpacket
	wire         video_in_decoder_avalon_decoder_source_valid;                                                               // Video_In_Decoder:stream_out_valid -> Video_RGB_Resampler:stream_in_valid
	wire         video_in_decoder_avalon_decoder_source_startofpacket;                                                       // Video_In_Decoder:stream_out_startofpacket -> Video_RGB_Resampler:stream_in_startofpacket
	wire   [7:0] video_in_decoder_avalon_decoder_source_data;                                                                // Video_In_Decoder:stream_out_data -> Video_RGB_Resampler:stream_in_data
	wire         video_in_decoder_avalon_decoder_source_ready;                                                               // Video_RGB_Resampler:stream_in_ready -> Video_In_Decoder:stream_out_ready
	wire         cpu_instruction_master_waitrequest;                                                                         // CPU_instruction_master_translator:av_waitrequest -> CPU:i_waitrequest
	wire  [21:0] cpu_instruction_master_address;                                                                             // CPU:i_address -> CPU_instruction_master_translator:av_address
	wire         cpu_instruction_master_read;                                                                                // CPU:i_read -> CPU_instruction_master_translator:av_read
	wire  [31:0] cpu_instruction_master_readdata;                                                                            // CPU_instruction_master_translator:av_readdata -> CPU:i_readdata
	wire         cpu_data_master_waitrequest;                                                                                // CPU_data_master_translator:av_waitrequest -> CPU:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                                                                  // CPU:d_writedata -> CPU_data_master_translator:av_writedata
	wire  [21:0] cpu_data_master_address;                                                                                    // CPU:d_address -> CPU_data_master_translator:av_address
	wire         cpu_data_master_write;                                                                                      // CPU:d_write -> CPU_data_master_translator:av_write
	wire         cpu_data_master_read;                                                                                       // CPU:d_read -> CPU_data_master_translator:av_read
	wire  [31:0] cpu_data_master_readdata;                                                                                   // CPU_data_master_translator:av_readdata -> CPU:d_readdata
	wire         cpu_data_master_debugaccess;                                                                                // CPU:jtag_debug_module_debugaccess_to_roms -> CPU_data_master_translator:av_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                                                                 // CPU:d_byteenable -> CPU_data_master_translator:av_byteenable
	wire         pixel_buffer_dma_avalon_pixel_dma_master_waitrequest;                                                       // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:av_waitrequest -> Pixel_Buffer_DMA:master_waitrequest
	wire  [31:0] pixel_buffer_dma_avalon_pixel_dma_master_address;                                                           // Pixel_Buffer_DMA:master_address -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:av_address
	wire         pixel_buffer_dma_avalon_pixel_dma_master_lock;                                                              // Pixel_Buffer_DMA:master_arbiterlock -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:av_lock
	wire         pixel_buffer_dma_avalon_pixel_dma_master_read;                                                              // Pixel_Buffer_DMA:master_read -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:av_read
	wire  [15:0] pixel_buffer_dma_avalon_pixel_dma_master_readdata;                                                          // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:av_readdata -> Pixel_Buffer_DMA:master_readdata
	wire         pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid;                                                     // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:av_readdatavalid -> Pixel_Buffer_DMA:master_readdatavalid
	wire         video_dma_avalon_dma_master_waitrequest;                                                                    // Video_DMA_avalon_dma_master_translator:av_waitrequest -> Video_DMA:master_waitrequest
	wire  [15:0] video_dma_avalon_dma_master_writedata;                                                                      // Video_DMA:master_writedata -> Video_DMA_avalon_dma_master_translator:av_writedata
	wire  [31:0] video_dma_avalon_dma_master_address;                                                                        // Video_DMA:master_address -> Video_DMA_avalon_dma_master_translator:av_address
	wire         video_dma_avalon_dma_master_write;                                                                          // Video_DMA:master_write -> Video_DMA_avalon_dma_master_translator:av_write
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                             // CPU_jtag_debug_module_translator:av_writedata -> CPU:jtag_debug_module_writedata
	wire   [8:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                               // CPU_jtag_debug_module_translator:av_address -> CPU:jtag_debug_module_address
	wire         cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                            // CPU_jtag_debug_module_translator:av_chipselect -> CPU:jtag_debug_module_select
	wire         cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                                 // CPU_jtag_debug_module_translator:av_write -> CPU:jtag_debug_module_write
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                              // CPU:jtag_debug_module_readdata -> CPU_jtag_debug_module_translator:av_readdata
	wire         cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                         // CPU_jtag_debug_module_translator:av_begintransfer -> CPU:jtag_debug_module_begintransfer
	wire         cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                           // CPU_jtag_debug_module_translator:av_debugaccess -> CPU:jtag_debug_module_debugaccess
	wire   [3:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                            // CPU_jtag_debug_module_translator:av_byteenable -> CPU:jtag_debug_module_byteenable
	wire  [31:0] onchip_memory_s1_translator_avalon_anti_slave_0_writedata;                                                  // Onchip_Memory_s1_translator:av_writedata -> Onchip_Memory:writedata
	wire  [11:0] onchip_memory_s1_translator_avalon_anti_slave_0_address;                                                    // Onchip_Memory_s1_translator:av_address -> Onchip_Memory:address
	wire         onchip_memory_s1_translator_avalon_anti_slave_0_chipselect;                                                 // Onchip_Memory_s1_translator:av_chipselect -> Onchip_Memory:chipselect
	wire         onchip_memory_s1_translator_avalon_anti_slave_0_clken;                                                      // Onchip_Memory_s1_translator:av_clken -> Onchip_Memory:clken
	wire         onchip_memory_s1_translator_avalon_anti_slave_0_write;                                                      // Onchip_Memory_s1_translator:av_write -> Onchip_Memory:write
	wire  [31:0] onchip_memory_s1_translator_avalon_anti_slave_0_readdata;                                                   // Onchip_Memory:readdata -> Onchip_Memory_s1_translator:av_readdata
	wire   [3:0] onchip_memory_s1_translator_avalon_anti_slave_0_byteenable;                                                 // Onchip_Memory_s1_translator:av_byteenable -> Onchip_Memory:byteenable
	wire  [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata;                                    // Pixel_Buffer_avalon_sram_slave_translator:av_writedata -> Pixel_Buffer:writedata
	wire  [19:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address;                                      // Pixel_Buffer_avalon_sram_slave_translator:av_address -> Pixel_Buffer:address
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write;                                        // Pixel_Buffer_avalon_sram_slave_translator:av_write -> Pixel_Buffer:write
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read;                                         // Pixel_Buffer_avalon_sram_slave_translator:av_read -> Pixel_Buffer:read
	wire  [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata;                                     // Pixel_Buffer:readdata -> Pixel_Buffer_avalon_sram_slave_translator:av_readdata
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid;                                // Pixel_Buffer:readdatavalid -> Pixel_Buffer_avalon_sram_slave_translator:av_readdatavalid
	wire   [1:0] pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable;                                   // Pixel_Buffer_avalon_sram_slave_translator:av_byteenable -> Pixel_Buffer:byteenable
	wire         av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest;                                // AV_Config:waitrequest -> AV_Config_avalon_av_config_slave_translator:av_waitrequest
	wire  [31:0] av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata;                                  // AV_Config_avalon_av_config_slave_translator:av_writedata -> AV_Config:writedata
	wire   [1:0] av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_address;                                    // AV_Config_avalon_av_config_slave_translator:av_address -> AV_Config:address
	wire         av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_write;                                      // AV_Config_avalon_av_config_slave_translator:av_write -> AV_Config:write
	wire         av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_read;                                       // AV_Config_avalon_av_config_slave_translator:av_read -> AV_Config:read
	wire  [31:0] av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata;                                   // AV_Config:readdata -> AV_Config_avalon_av_config_slave_translator:av_readdata
	wire   [3:0] av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable;                                 // AV_Config_avalon_av_config_slave_translator:av_byteenable -> AV_Config:byteenable
	wire  [31:0] video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata;                                // Video_DMA_avalon_dma_control_slave_translator:av_writedata -> Video_DMA:slave_writedata
	wire   [1:0] video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_address;                                  // Video_DMA_avalon_dma_control_slave_translator:av_address -> Video_DMA:slave_address
	wire         video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_write;                                    // Video_DMA_avalon_dma_control_slave_translator:av_write -> Video_DMA:slave_write
	wire         video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_read;                                     // Video_DMA_avalon_dma_control_slave_translator:av_read -> Video_DMA:slave_read
	wire  [31:0] video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata;                                 // Video_DMA:slave_readdata -> Video_DMA_avalon_dma_control_slave_translator:av_readdata
	wire   [3:0] video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable;                               // Video_DMA_avalon_dma_control_slave_translator:av_byteenable -> Video_DMA:slave_byteenable
	wire  [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_writedata;                             // Pixel_Buffer_DMA_avalon_control_slave_translator:av_writedata -> Pixel_Buffer_DMA:slave_writedata
	wire   [1:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_address;                               // Pixel_Buffer_DMA_avalon_control_slave_translator:av_address -> Pixel_Buffer_DMA:slave_address
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_write;                                 // Pixel_Buffer_DMA_avalon_control_slave_translator:av_write -> Pixel_Buffer_DMA:slave_write
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_read;                                  // Pixel_Buffer_DMA_avalon_control_slave_translator:av_read -> Pixel_Buffer_DMA:slave_read
	wire  [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_readdata;                              // Pixel_Buffer_DMA:slave_readdata -> Pixel_Buffer_DMA_avalon_control_slave_translator:av_readdata
	wire   [3:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_byteenable;                            // Pixel_Buffer_DMA_avalon_control_slave_translator:av_byteenable -> Pixel_Buffer_DMA:slave_byteenable
	wire         cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                                    // CPU_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> CPU_instruction_master_translator:uav_waitrequest
	wire   [2:0] cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                                     // CPU_instruction_master_translator:uav_burstcount -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_instruction_master_translator_avalon_universal_master_0_writedata;                                      // CPU_instruction_master_translator:uav_writedata -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] cpu_instruction_master_translator_avalon_universal_master_0_address;                                        // CPU_instruction_master_translator:uav_address -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_instruction_master_translator_avalon_universal_master_0_lock;                                           // CPU_instruction_master_translator:uav_lock -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_instruction_master_translator_avalon_universal_master_0_write;                                          // CPU_instruction_master_translator:uav_write -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_instruction_master_translator_avalon_universal_master_0_read;                                           // CPU_instruction_master_translator:uav_read -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_instruction_master_translator_avalon_universal_master_0_readdata;                                       // CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> CPU_instruction_master_translator:uav_readdata
	wire         cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                                    // CPU_instruction_master_translator:uav_debugaccess -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                                     // CPU_instruction_master_translator:uav_byteenable -> CPU_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                                  // CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> CPU_instruction_master_translator:uav_readdatavalid
	wire         cpu_data_master_translator_avalon_universal_master_0_waitrequest;                                           // CPU_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> CPU_data_master_translator:uav_waitrequest
	wire   [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                                            // CPU_data_master_translator:uav_burstcount -> CPU_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                                             // CPU_data_master_translator:uav_writedata -> CPU_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] cpu_data_master_translator_avalon_universal_master_0_address;                                               // CPU_data_master_translator:uav_address -> CPU_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_data_master_translator_avalon_universal_master_0_lock;                                                  // CPU_data_master_translator:uav_lock -> CPU_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_data_master_translator_avalon_universal_master_0_write;                                                 // CPU_data_master_translator:uav_write -> CPU_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_data_master_translator_avalon_universal_master_0_read;                                                  // CPU_data_master_translator:uav_read -> CPU_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                                              // CPU_data_master_translator_avalon_universal_master_0_agent:av_readdata -> CPU_data_master_translator:uav_readdata
	wire         cpu_data_master_translator_avalon_universal_master_0_debugaccess;                                           // CPU_data_master_translator:uav_debugaccess -> CPU_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                                            // CPU_data_master_translator:uav_byteenable -> CPU_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                                         // CPU_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> CPU_data_master_translator:uav_readdatavalid
	wire         pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest;                  // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_waitrequest
	wire   [1:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount;                   // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_burstcount -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [15:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata;                    // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_writedata -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address;                      // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_address -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire         pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock;                         // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_lock -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire         pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write;                        // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_write -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire         pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read;                         // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_read -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire  [15:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata;                     // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_readdata
	wire         pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess;                  // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_debugaccess -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [1:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable;                   // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_byteenable -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid;                // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:uav_readdatavalid
	wire         video_dma_avalon_dma_master_translator_avalon_universal_master_0_waitrequest;                               // Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_waitrequest -> Video_DMA_avalon_dma_master_translator:uav_waitrequest
	wire   [1:0] video_dma_avalon_dma_master_translator_avalon_universal_master_0_burstcount;                                // Video_DMA_avalon_dma_master_translator:uav_burstcount -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [15:0] video_dma_avalon_dma_master_translator_avalon_universal_master_0_writedata;                                 // Video_DMA_avalon_dma_master_translator:uav_writedata -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] video_dma_avalon_dma_master_translator_avalon_universal_master_0_address;                                   // Video_DMA_avalon_dma_master_translator:uav_address -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_address
	wire         video_dma_avalon_dma_master_translator_avalon_universal_master_0_lock;                                      // Video_DMA_avalon_dma_master_translator:uav_lock -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_lock
	wire         video_dma_avalon_dma_master_translator_avalon_universal_master_0_write;                                     // Video_DMA_avalon_dma_master_translator:uav_write -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_write
	wire         video_dma_avalon_dma_master_translator_avalon_universal_master_0_read;                                      // Video_DMA_avalon_dma_master_translator:uav_read -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_read
	wire  [15:0] video_dma_avalon_dma_master_translator_avalon_universal_master_0_readdata;                                  // Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdata -> Video_DMA_avalon_dma_master_translator:uav_readdata
	wire         video_dma_avalon_dma_master_translator_avalon_universal_master_0_debugaccess;                               // Video_DMA_avalon_dma_master_translator:uav_debugaccess -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [1:0] video_dma_avalon_dma_master_translator_avalon_universal_master_0_byteenable;                                // Video_DMA_avalon_dma_master_translator:uav_byteenable -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         video_dma_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid;                             // Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> Video_DMA_avalon_dma_master_translator:uav_readdatavalid
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // CPU_jtag_debug_module_translator:uav_waitrequest -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> CPU_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                               // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> CPU_jtag_debug_module_translator:uav_writedata
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                                 // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> CPU_jtag_debug_module_translator:uav_address
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                   // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> CPU_jtag_debug_module_translator:uav_write
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                    // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> CPU_jtag_debug_module_translator:uav_lock
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                    // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> CPU_jtag_debug_module_translator:uav_read
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                                // CPU_jtag_debug_module_translator:uav_readdata -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // CPU_jtag_debug_module_translator:uav_readdatavalid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CPU_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> CPU_jtag_debug_module_translator:uav_byteenable
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                             // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // Onchip_Memory_s1_translator:uav_waitrequest -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> Onchip_Memory_s1_translator:uav_burstcount
	wire  [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> Onchip_Memory_s1_translator:uav_writedata
	wire  [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> Onchip_Memory_s1_translator:uav_address
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> Onchip_Memory_s1_translator:uav_write
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> Onchip_Memory_s1_translator:uav_lock
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> Onchip_Memory_s1_translator:uav_read
	wire  [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // Onchip_Memory_s1_translator:uav_readdata -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // Onchip_Memory_s1_translator:uav_readdatavalid -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Onchip_Memory_s1_translator:uav_debugaccess
	wire   [3:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> Onchip_Memory_s1_translator:uav_byteenable
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // Pixel_Buffer_avalon_sram_slave_translator:uav_waitrequest -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Pixel_Buffer_avalon_sram_slave_translator:uav_burstcount
	wire  [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                      // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Pixel_Buffer_avalon_sram_slave_translator:uav_writedata
	wire  [31:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address;                        // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_address -> Pixel_Buffer_avalon_sram_slave_translator:uav_address
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write;                          // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_write -> Pixel_Buffer_avalon_sram_slave_translator:uav_write
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock;                           // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Pixel_Buffer_avalon_sram_slave_translator:uav_lock
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read;                           // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_read -> Pixel_Buffer_avalon_sram_slave_translator:uav_read
	wire  [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                       // Pixel_Buffer_avalon_sram_slave_translator:uav_readdata -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // Pixel_Buffer_avalon_sram_slave_translator:uav_readdatavalid -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Pixel_Buffer_avalon_sram_slave_translator:uav_debugaccess
	wire   [1:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Pixel_Buffer_avalon_sram_slave_translator:uav_byteenable
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [69:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                    // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [69:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [15:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // AV_Config_avalon_av_config_slave_translator:uav_waitrequest -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> AV_Config_avalon_av_config_slave_translator:uav_burstcount
	wire  [31:0] av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                    // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> AV_Config_avalon_av_config_slave_translator:uav_writedata
	wire  [31:0] av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address;                      // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_address -> AV_Config_avalon_av_config_slave_translator:uav_address
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write;                        // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_write -> AV_Config_avalon_av_config_slave_translator:uav_write
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock;                         // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_lock -> AV_Config_avalon_av_config_slave_translator:uav_lock
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read;                         // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_read -> AV_Config_avalon_av_config_slave_translator:uav_read
	wire  [31:0] av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                     // AV_Config_avalon_av_config_slave_translator:uav_readdata -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // AV_Config_avalon_av_config_slave_translator:uav_readdatavalid -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> AV_Config_avalon_av_config_slave_translator:uav_debugaccess
	wire   [3:0] av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> AV_Config_avalon_av_config_slave_translator:uav_byteenable
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                  // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // Video_DMA_avalon_dma_control_slave_translator:uav_waitrequest -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Video_DMA_avalon_dma_control_slave_translator:uav_burstcount
	wire  [31:0] video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                  // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Video_DMA_avalon_dma_control_slave_translator:uav_writedata
	wire  [31:0] video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                    // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> Video_DMA_avalon_dma_control_slave_translator:uav_address
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                      // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> Video_DMA_avalon_dma_control_slave_translator:uav_write
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                       // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Video_DMA_avalon_dma_control_slave_translator:uav_lock
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                       // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> Video_DMA_avalon_dma_control_slave_translator:uav_read
	wire  [31:0] video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                   // Video_DMA_avalon_dma_control_slave_translator:uav_readdata -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // Video_DMA_avalon_dma_control_slave_translator:uav_readdatavalid -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Video_DMA_avalon_dma_control_slave_translator:uav_debugaccess
	wire   [3:0] video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Video_DMA_avalon_dma_control_slave_translator:uav_byteenable
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;               // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;               // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Pixel_Buffer_DMA_avalon_control_slave_translator:uav_waitrequest -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_burstcount
	wire  [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_writedata
	wire  [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_address
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_write
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_lock
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_read
	wire  [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // Pixel_Buffer_DMA_avalon_control_slave_translator:uav_readdata -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Pixel_Buffer_DMA_avalon_control_slave_translator:uav_readdatavalid -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_debugaccess
	wire   [3:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Pixel_Buffer_DMA_avalon_control_slave_translator:uav_byteenable
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                           // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                                 // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                         // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [86:0] cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                                  // CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                                 // addr_router:sink_ready -> CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                  // CPU_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                        // CPU_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                // CPU_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [86:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                                         // CPU_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                        // addr_router_001:sink_ready -> CPU_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;         // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire         pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid;               // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire         pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket;       // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [68:0] pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data;                // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire         pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready;               // addr_router_002:sink_ready -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire         video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid;                            // Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire         video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [68:0] video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data;                             // Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire         video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router_003:sink_ready -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                   // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [86:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                    // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router:sink_ready -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [86:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_001:sink_ready -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid;                          // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [68:0] pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data;                           // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_002:sink_ready -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid;                        // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [86:0] av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data;                         // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready;                        // id_router_003:sink_ready -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                      // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [86:0] video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                       // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_004:sink_ready -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [86:0] pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_005:sink_ready -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                                // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                                      // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                              // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [86:0] addr_router_src_data;                                                                                       // addr_router:src_data -> limiter:cmd_sink_data
	wire   [5:0] addr_router_src_channel;                                                                                    // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                                      // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                                // limiter:rsp_src_endofpacket -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                                      // limiter:rsp_src_valid -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                              // limiter:rsp_src_startofpacket -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [86:0] limiter_rsp_src_data;                                                                                       // limiter:rsp_src_data -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [5:0] limiter_rsp_src_channel;                                                                                    // limiter:rsp_src_channel -> CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                                      // CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         addr_router_001_src_endofpacket;                                                                            // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire         addr_router_001_src_valid;                                                                                  // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire         addr_router_001_src_startofpacket;                                                                          // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [86:0] addr_router_001_src_data;                                                                                   // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire   [5:0] addr_router_001_src_channel;                                                                                // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire         addr_router_001_src_ready;                                                                                  // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire         limiter_001_rsp_src_endofpacket;                                                                            // limiter_001:rsp_src_endofpacket -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_001_rsp_src_valid;                                                                                  // limiter_001:rsp_src_valid -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_001_rsp_src_startofpacket;                                                                          // limiter_001:rsp_src_startofpacket -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [86:0] limiter_001_rsp_src_data;                                                                                   // limiter_001:rsp_src_data -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [5:0] limiter_001_rsp_src_channel;                                                                                // limiter_001:rsp_src_channel -> CPU_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_001_rsp_src_ready;                                                                                  // CPU_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire         addr_router_002_src_endofpacket;                                                                            // addr_router_002:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	wire         addr_router_002_src_valid;                                                                                  // addr_router_002:src_valid -> limiter_002:cmd_sink_valid
	wire         addr_router_002_src_startofpacket;                                                                          // addr_router_002:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	wire  [68:0] addr_router_002_src_data;                                                                                   // addr_router_002:src_data -> limiter_002:cmd_sink_data
	wire   [5:0] addr_router_002_src_channel;                                                                                // addr_router_002:src_channel -> limiter_002:cmd_sink_channel
	wire         addr_router_002_src_ready;                                                                                  // limiter_002:cmd_sink_ready -> addr_router_002:src_ready
	wire         limiter_002_rsp_src_endofpacket;                                                                            // limiter_002:rsp_src_endofpacket -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_002_rsp_src_valid;                                                                                  // limiter_002:rsp_src_valid -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_002_rsp_src_startofpacket;                                                                          // limiter_002:rsp_src_startofpacket -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [68:0] limiter_002_rsp_src_data;                                                                                   // limiter_002:rsp_src_data -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [5:0] limiter_002_rsp_src_channel;                                                                                // limiter_002:rsp_src_channel -> Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_002_rsp_src_ready;                                                                                  // Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_002:rsp_src_ready
	wire         addr_router_003_src_endofpacket;                                                                            // addr_router_003:src_endofpacket -> limiter_003:cmd_sink_endofpacket
	wire         addr_router_003_src_valid;                                                                                  // addr_router_003:src_valid -> limiter_003:cmd_sink_valid
	wire         addr_router_003_src_startofpacket;                                                                          // addr_router_003:src_startofpacket -> limiter_003:cmd_sink_startofpacket
	wire  [68:0] addr_router_003_src_data;                                                                                   // addr_router_003:src_data -> limiter_003:cmd_sink_data
	wire   [5:0] addr_router_003_src_channel;                                                                                // addr_router_003:src_channel -> limiter_003:cmd_sink_channel
	wire         addr_router_003_src_ready;                                                                                  // limiter_003:cmd_sink_ready -> addr_router_003:src_ready
	wire         limiter_003_rsp_src_endofpacket;                                                                            // limiter_003:rsp_src_endofpacket -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_003_rsp_src_valid;                                                                                  // limiter_003:rsp_src_valid -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_003_rsp_src_startofpacket;                                                                          // limiter_003:rsp_src_startofpacket -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [68:0] limiter_003_rsp_src_data;                                                                                   // limiter_003:rsp_src_data -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [5:0] limiter_003_rsp_src_channel;                                                                                // limiter_003:rsp_src_channel -> Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_003_rsp_src_ready;                                                                                  // Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_003:rsp_src_ready
	wire         burst_adapter_source0_endofpacket;                                                                          // burst_adapter:source0_endofpacket -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_source0_valid;                                                                                // burst_adapter:source0_valid -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_source0_startofpacket;                                                                        // burst_adapter:source0_startofpacket -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [68:0] burst_adapter_source0_data;                                                                                 // burst_adapter:source0_data -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_source0_ready;                                                                                // Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [5:0] burst_adapter_source0_channel;                                                                              // burst_adapter:source0_channel -> Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rst_controller_reset_out_reset;                                                                             // rst_controller:reset_out -> [AV_Config:reset, AV_Config_avalon_av_config_slave_translator:reset, AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:reset, AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CPU:reset_n, CPU_data_master_translator:reset, CPU_data_master_translator_avalon_universal_master_0_agent:reset, CPU_instruction_master_translator:reset, CPU_instruction_master_translator_avalon_universal_master_0_agent:reset, CPU_jtag_debug_module_translator:reset, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Dual_Clock_FIFO:reset_stream_in, Onchip_Memory:reset, Onchip_Memory_s1_translator:reset, Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:reset, Onchip_Memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Pixel_Buffer:reset, Pixel_Buffer_DMA:reset, Pixel_Buffer_DMA_avalon_control_slave_translator:reset, Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:reset, Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Pixel_Buffer_DMA_avalon_pixel_dma_master_translator:reset, Pixel_Buffer_DMA_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent:reset, Pixel_Buffer_avalon_sram_slave_translator:reset, Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent:reset, Pixel_Buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Pixel_RGB_Resampler:reset, Pixel_Scaler:reset, Video_Clipper:reset, Video_DMA:reset, Video_DMA_avalon_dma_control_slave_translator:reset, Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:reset, Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Video_DMA_avalon_dma_master_translator:reset, Video_DMA_avalon_dma_master_translator_avalon_universal_master_0_agent:reset, Video_In_Decoder:reset, Video_RGB_Resampler:reset, Video_Scaler:reset, addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, irq_mapper:reset, limiter:reset, limiter_001:reset, limiter_002:reset, limiter_003:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, width_adapter:reset, width_adapter_001:reset]
	wire         cpu_jtag_debug_module_reset_reset;                                                                          // CPU:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	wire         rst_controller_001_reset_out_reset;                                                                         // rst_controller_001:reset_out -> [Dual_Clock_FIFO:reset_stream_out, VGA_Controller:reset]
	wire         rst_controller_002_reset_out_reset;                                                                         // rst_controller_002:reset_out -> Clock_Signals:reset
	wire         cmd_xbar_demux_src0_endofpacket;                                                                            // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                                  // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                          // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [86:0] cmd_xbar_demux_src0_data;                                                                                   // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [5:0] cmd_xbar_demux_src0_channel;                                                                                // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                                  // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                            // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                                  // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                          // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [86:0] cmd_xbar_demux_src1_data;                                                                                   // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [5:0] cmd_xbar_demux_src1_channel;                                                                                // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                                  // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                        // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                              // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                                      // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [86:0] cmd_xbar_demux_001_src0_data;                                                                               // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [5:0] cmd_xbar_demux_001_src0_channel;                                                                            // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                              // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                        // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                              // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                                      // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [86:0] cmd_xbar_demux_001_src1_data;                                                                               // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [5:0] cmd_xbar_demux_001_src1_channel;                                                                            // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                              // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                        // cmd_xbar_demux_001:src3_endofpacket -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                              // cmd_xbar_demux_001:src3_valid -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                                      // cmd_xbar_demux_001:src3_startofpacket -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_001_src3_data;                                                                               // cmd_xbar_demux_001:src3_data -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] cmd_xbar_demux_001_src3_channel;                                                                            // cmd_xbar_demux_001:src3_channel -> AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                        // cmd_xbar_demux_001:src4_endofpacket -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                              // cmd_xbar_demux_001:src4_valid -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                                      // cmd_xbar_demux_001:src4_startofpacket -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_001_src4_data;                                                                               // cmd_xbar_demux_001:src4_data -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] cmd_xbar_demux_001_src4_channel;                                                                            // cmd_xbar_demux_001:src4_channel -> Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                        // cmd_xbar_demux_001:src5_endofpacket -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                              // cmd_xbar_demux_001:src5_valid -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                                      // cmd_xbar_demux_001:src5_startofpacket -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_001_src5_data;                                                                               // cmd_xbar_demux_001:src5_data -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] cmd_xbar_demux_001_src5_channel;                                                                            // cmd_xbar_demux_001:src5_channel -> Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_002_src0_endofpacket;                                                                        // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_002_src0_valid;                                                                              // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_002_src0_startofpacket;                                                                      // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [68:0] cmd_xbar_demux_002_src0_data;                                                                               // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_002:sink1_data
	wire   [5:0] cmd_xbar_demux_002_src0_channel;                                                                            // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_002_src0_ready;                                                                              // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire         cmd_xbar_demux_003_src0_endofpacket;                                                                        // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_002:sink2_endofpacket
	wire         cmd_xbar_demux_003_src0_valid;                                                                              // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_002:sink2_valid
	wire         cmd_xbar_demux_003_src0_startofpacket;                                                                      // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_002:sink2_startofpacket
	wire  [68:0] cmd_xbar_demux_003_src0_data;                                                                               // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_002:sink2_data
	wire   [5:0] cmd_xbar_demux_003_src0_channel;                                                                            // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_002:sink2_channel
	wire         cmd_xbar_demux_003_src0_ready;                                                                              // cmd_xbar_mux_002:sink2_ready -> cmd_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_src0_endofpacket;                                                                            // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                                  // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                          // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [86:0] rsp_xbar_demux_src0_data;                                                                                   // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [5:0] rsp_xbar_demux_src0_channel;                                                                                // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                                  // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                            // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                                  // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                          // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [86:0] rsp_xbar_demux_src1_data;                                                                                   // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [5:0] rsp_xbar_demux_src1_channel;                                                                                // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                                  // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                        // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                              // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                                      // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [86:0] rsp_xbar_demux_001_src0_data;                                                                               // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [5:0] rsp_xbar_demux_001_src0_channel;                                                                            // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                              // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                        // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                              // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                                      // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [86:0] rsp_xbar_demux_001_src1_data;                                                                               // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [5:0] rsp_xbar_demux_001_src1_channel;                                                                            // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                              // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                                        // rsp_xbar_demux_002:src1_endofpacket -> limiter_002:rsp_sink_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                              // rsp_xbar_demux_002:src1_valid -> limiter_002:rsp_sink_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                                      // rsp_xbar_demux_002:src1_startofpacket -> limiter_002:rsp_sink_startofpacket
	wire  [68:0] rsp_xbar_demux_002_src1_data;                                                                               // rsp_xbar_demux_002:src1_data -> limiter_002:rsp_sink_data
	wire   [5:0] rsp_xbar_demux_002_src1_channel;                                                                            // rsp_xbar_demux_002:src1_channel -> limiter_002:rsp_sink_channel
	wire         rsp_xbar_demux_002_src2_endofpacket;                                                                        // rsp_xbar_demux_002:src2_endofpacket -> limiter_003:rsp_sink_endofpacket
	wire         rsp_xbar_demux_002_src2_valid;                                                                              // rsp_xbar_demux_002:src2_valid -> limiter_003:rsp_sink_valid
	wire         rsp_xbar_demux_002_src2_startofpacket;                                                                      // rsp_xbar_demux_002:src2_startofpacket -> limiter_003:rsp_sink_startofpacket
	wire  [68:0] rsp_xbar_demux_002_src2_data;                                                                               // rsp_xbar_demux_002:src2_data -> limiter_003:rsp_sink_data
	wire   [5:0] rsp_xbar_demux_002_src2_channel;                                                                            // rsp_xbar_demux_002:src2_channel -> limiter_003:rsp_sink_channel
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                        // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                              // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                                      // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [86:0] rsp_xbar_demux_003_src0_data;                                                                               // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [5:0] rsp_xbar_demux_003_src0_channel;                                                                            // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                              // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                        // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                              // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                                      // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [86:0] rsp_xbar_demux_004_src0_data;                                                                               // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [5:0] rsp_xbar_demux_004_src0_channel;                                                                            // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                              // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                        // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                              // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                                      // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [86:0] rsp_xbar_demux_005_src0_data;                                                                               // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [5:0] rsp_xbar_demux_005_src0_channel;                                                                            // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                              // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                                // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                              // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [86:0] limiter_cmd_src_data;                                                                                       // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [5:0] limiter_cmd_src_channel;                                                                                    // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                                      // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                               // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                                     // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                             // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [86:0] rsp_xbar_mux_src_data;                                                                                      // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [5:0] rsp_xbar_mux_src_channel;                                                                                   // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                                     // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         limiter_001_cmd_src_endofpacket;                                                                            // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         limiter_001_cmd_src_startofpacket;                                                                          // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [86:0] limiter_001_cmd_src_data;                                                                                   // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire   [5:0] limiter_001_cmd_src_channel;                                                                                // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire         limiter_001_cmd_src_ready;                                                                                  // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                           // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                                 // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                         // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [86:0] rsp_xbar_mux_001_src_data;                                                                                  // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire   [5:0] rsp_xbar_mux_001_src_channel;                                                                               // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                                 // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire         limiter_002_cmd_src_endofpacket;                                                                            // limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire         limiter_002_cmd_src_startofpacket;                                                                          // limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [68:0] limiter_002_cmd_src_data;                                                                                   // limiter_002:cmd_src_data -> cmd_xbar_demux_002:sink_data
	wire   [5:0] limiter_002_cmd_src_channel;                                                                                // limiter_002:cmd_src_channel -> cmd_xbar_demux_002:sink_channel
	wire         limiter_002_cmd_src_ready;                                                                                  // cmd_xbar_demux_002:sink_ready -> limiter_002:cmd_src_ready
	wire         rsp_xbar_demux_002_src1_ready;                                                                              // limiter_002:rsp_sink_ready -> rsp_xbar_demux_002:src1_ready
	wire         limiter_003_cmd_src_endofpacket;                                                                            // limiter_003:cmd_src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire         limiter_003_cmd_src_startofpacket;                                                                          // limiter_003:cmd_src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [68:0] limiter_003_cmd_src_data;                                                                                   // limiter_003:cmd_src_data -> cmd_xbar_demux_003:sink_data
	wire   [5:0] limiter_003_cmd_src_channel;                                                                                // limiter_003:cmd_src_channel -> cmd_xbar_demux_003:sink_channel
	wire         limiter_003_cmd_src_ready;                                                                                  // cmd_xbar_demux_003:sink_ready -> limiter_003:cmd_src_ready
	wire         rsp_xbar_demux_002_src2_ready;                                                                              // limiter_003:rsp_sink_ready -> rsp_xbar_demux_002:src2_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                               // cmd_xbar_mux:src_endofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                                     // cmd_xbar_mux:src_valid -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                             // cmd_xbar_mux:src_startofpacket -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_mux_src_data;                                                                                      // cmd_xbar_mux:src_data -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] cmd_xbar_mux_src_channel;                                                                                   // cmd_xbar_mux:src_channel -> CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                                     // CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                                  // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                        // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                                // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [86:0] id_router_src_data;                                                                                         // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [5:0] id_router_src_channel;                                                                                      // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                        // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                           // cmd_xbar_mux_001:src_endofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                                 // cmd_xbar_mux_001:src_valid -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                         // cmd_xbar_mux_001:src_startofpacket -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_mux_001_src_data;                                                                                  // cmd_xbar_mux_001:src_data -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] cmd_xbar_mux_001_src_channel;                                                                               // cmd_xbar_mux_001:src_channel -> Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                                 // Onchip_Memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                              // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                                    // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                            // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [86:0] id_router_001_src_data;                                                                                     // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [5:0] id_router_001_src_channel;                                                                                  // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                                    // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                           // cmd_xbar_mux_002:src_endofpacket -> burst_adapter:sink0_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                                 // cmd_xbar_mux_002:src_valid -> burst_adapter:sink0_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                         // cmd_xbar_mux_002:src_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [68:0] cmd_xbar_mux_002_src_data;                                                                                  // cmd_xbar_mux_002:src_data -> burst_adapter:sink0_data
	wire   [5:0] cmd_xbar_mux_002_src_channel;                                                                               // cmd_xbar_mux_002:src_channel -> burst_adapter:sink0_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                                 // burst_adapter:sink0_ready -> cmd_xbar_mux_002:src_ready
	wire         id_router_002_src_endofpacket;                                                                              // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                                    // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                            // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [68:0] id_router_002_src_data;                                                                                     // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [5:0] id_router_002_src_channel;                                                                                  // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                                    // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_001_src3_ready;                                                                              // AV_Config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire         id_router_003_src_endofpacket;                                                                              // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                                    // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                            // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [86:0] id_router_003_src_data;                                                                                     // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [5:0] id_router_003_src_channel;                                                                                  // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                                    // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_001_src4_ready;                                                                              // Video_DMA_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire         id_router_004_src_endofpacket;                                                                              // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                                    // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                            // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [86:0] id_router_004_src_data;                                                                                     // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [5:0] id_router_004_src_channel;                                                                                  // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                                    // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_001_src5_ready;                                                                              // Pixel_Buffer_DMA_avalon_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire         id_router_005_src_endofpacket;                                                                              // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                                    // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                            // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [86:0] id_router_005_src_data;                                                                                     // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [5:0] id_router_005_src_channel;                                                                                  // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                                    // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                        // cmd_xbar_demux_001:src2_endofpacket -> width_adapter:in_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                              // cmd_xbar_demux_001:src2_valid -> width_adapter:in_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                                      // cmd_xbar_demux_001:src2_startofpacket -> width_adapter:in_startofpacket
	wire  [86:0] cmd_xbar_demux_001_src2_data;                                                                               // cmd_xbar_demux_001:src2_data -> width_adapter:in_data
	wire   [5:0] cmd_xbar_demux_001_src2_channel;                                                                            // cmd_xbar_demux_001:src2_channel -> width_adapter:in_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                              // width_adapter:in_ready -> cmd_xbar_demux_001:src2_ready
	wire         width_adapter_src_endofpacket;                                                                              // width_adapter:out_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         width_adapter_src_valid;                                                                                    // width_adapter:out_valid -> cmd_xbar_mux_002:sink0_valid
	wire         width_adapter_src_startofpacket;                                                                            // width_adapter:out_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [68:0] width_adapter_src_data;                                                                                     // width_adapter:out_data -> cmd_xbar_mux_002:sink0_data
	wire         width_adapter_src_ready;                                                                                    // cmd_xbar_mux_002:sink0_ready -> width_adapter:out_ready
	wire   [5:0] width_adapter_src_channel;                                                                                  // width_adapter:out_channel -> cmd_xbar_mux_002:sink0_channel
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                        // rsp_xbar_demux_002:src0_endofpacket -> width_adapter_001:in_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                              // rsp_xbar_demux_002:src0_valid -> width_adapter_001:in_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                                      // rsp_xbar_demux_002:src0_startofpacket -> width_adapter_001:in_startofpacket
	wire  [68:0] rsp_xbar_demux_002_src0_data;                                                                               // rsp_xbar_demux_002:src0_data -> width_adapter_001:in_data
	wire   [5:0] rsp_xbar_demux_002_src0_channel;                                                                            // rsp_xbar_demux_002:src0_channel -> width_adapter_001:in_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                              // width_adapter_001:in_ready -> rsp_xbar_demux_002:src0_ready
	wire         width_adapter_001_src_endofpacket;                                                                          // width_adapter_001:out_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         width_adapter_001_src_valid;                                                                                // width_adapter_001:out_valid -> rsp_xbar_mux_001:sink2_valid
	wire         width_adapter_001_src_startofpacket;                                                                        // width_adapter_001:out_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [86:0] width_adapter_001_src_data;                                                                                 // width_adapter_001:out_data -> rsp_xbar_mux_001:sink2_data
	wire         width_adapter_001_src_ready;                                                                                // rsp_xbar_mux_001:sink2_ready -> width_adapter_001:out_ready
	wire   [5:0] width_adapter_001_src_channel;                                                                              // width_adapter_001:out_channel -> rsp_xbar_mux_001:sink2_channel
	wire   [5:0] limiter_cmd_valid_data;                                                                                     // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [5:0] limiter_001_cmd_valid_data;                                                                                 // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire   [5:0] limiter_002_cmd_valid_data;                                                                                 // limiter_002:cmd_src_valid -> cmd_xbar_demux_002:sink_valid
	wire   [5:0] limiter_003_cmd_valid_data;                                                                                 // limiter_003:cmd_src_valid -> cmd_xbar_demux_003:sink_valid
	wire  [31:0] cpu_d_irq_irq;                                                                                              // irq_mapper:sender_irq -> CPU:d_irq

	Video_System_Onchip_Memory onchip_memory (
		.clk        (clock_signals_sys_clk_clk),                                  //   clk1.clk
		.address    (onchip_memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (onchip_memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (onchip_memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (onchip_memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (onchip_memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (onchip_memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                              // reset1.reset
	);

	Video_System_Dual_Clock_FIFO dual_clock_fifo (
		.clk_stream_in            (clock_signals_sys_clk_clk),                             //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                        //   clock_stream_in_reset.reset
		.clk_stream_out           (clock_signals_vga_clk_clk),                             //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_001_reset_out_reset),                    //  clock_stream_out_reset.reset
		.stream_in_ready          (pixel_scaler_avalon_scaler_source_ready),               //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (pixel_scaler_avalon_scaler_source_startofpacket),       //                        .startofpacket
		.stream_in_endofpacket    (pixel_scaler_avalon_scaler_source_endofpacket),         //                        .endofpacket
		.stream_in_valid          (pixel_scaler_avalon_scaler_source_valid),               //                        .valid
		.stream_in_data           (pixel_scaler_avalon_scaler_source_data),                //                        .data
		.stream_out_ready         (dual_clock_fifo_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (dual_clock_fifo_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (dual_clock_fifo_avalon_dc_buffer_source_data)           //                        .data
	);

	Video_System_Pixel_Buffer pixel_buffer (
		.clk           (clock_signals_sys_clk_clk),                                                   //        clock_reset.clk
		.reset         (rst_controller_reset_out_reset),                                              //  clock_reset_reset.reset
		.SRAM_DQ       (SRAM_DQ_to_and_from_the_Pixel_Buffer),                                        // external_interface.export
		.SRAM_ADDR     (SRAM_ADDR_from_the_Pixel_Buffer),                                             //                   .export
		.SRAM_LB_N     (SRAM_LB_N_from_the_Pixel_Buffer),                                             //                   .export
		.SRAM_UB_N     (SRAM_UB_N_from_the_Pixel_Buffer),                                             //                   .export
		.SRAM_CE_N     (SRAM_CE_N_from_the_Pixel_Buffer),                                             //                   .export
		.SRAM_OE_N     (SRAM_OE_N_from_the_Pixel_Buffer),                                             //                   .export
		.SRAM_WE_N     (SRAM_WE_N_from_the_Pixel_Buffer),                                             //                   .export
		.address       (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address),       //  avalon_sram_slave.address
		.byteenable    (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.read          (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read),          //                   .read
		.write         (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write),         //                   .write
		.writedata     (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.readdata      (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.readdatavalid (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid)  //                   .readdatavalid
	);

	Video_System_Pixel_Buffer_DMA pixel_buffer_dma (
		.clk                  (clock_signals_sys_clk_clk),                                                       //             clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                                                  //       clock_reset_reset.reset
		.master_readdatavalid (pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),                          // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),                            //                        .waitrequest
		.master_address       (pixel_buffer_dma_avalon_pixel_dma_master_address),                                //                        .address
		.master_arbiterlock   (pixel_buffer_dma_avalon_pixel_dma_master_lock),                                   //                        .lock
		.master_read          (pixel_buffer_dma_avalon_pixel_dma_master_read),                                   //                        .read
		.master_readdata      (pixel_buffer_dma_avalon_pixel_dma_master_readdata),                               //                        .readdata
		.slave_address        (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_address),    //    avalon_control_slave.address
		.slave_byteenable     (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_byteenable), //                        .byteenable
		.slave_read           (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_read),       //                        .read
		.slave_write          (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_write),      //                        .write
		.slave_writedata      (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_writedata),  //                        .writedata
		.slave_readdata       (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_readdata),   //                        .readdata
		.stream_ready         (pixel_buffer_dma_avalon_pixel_source_ready),                                      //     avalon_pixel_source.ready
		.stream_startofpacket (pixel_buffer_dma_avalon_pixel_source_startofpacket),                              //                        .startofpacket
		.stream_endofpacket   (pixel_buffer_dma_avalon_pixel_source_endofpacket),                                //                        .endofpacket
		.stream_valid         (pixel_buffer_dma_avalon_pixel_source_valid),                                      //                        .valid
		.stream_data          (pixel_buffer_dma_avalon_pixel_source_data)                                        //                        .data
	);

	Video_System_Pixel_RGB_Resampler pixel_rgb_resampler (
		.clk                      (clock_signals_sys_clk_clk),                           //       clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                      // clock_reset_reset.reset
		.stream_in_startofpacket  (pixel_buffer_dma_avalon_pixel_source_startofpacket),  //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (pixel_buffer_dma_avalon_pixel_source_endofpacket),    //                  .endofpacket
		.stream_in_valid          (pixel_buffer_dma_avalon_pixel_source_valid),          //                  .valid
		.stream_in_ready          (pixel_buffer_dma_avalon_pixel_source_ready),          //                  .ready
		.stream_in_data           (pixel_buffer_dma_avalon_pixel_source_data),           //                  .data
		.stream_out_ready         (pixel_rgb_resampler_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (pixel_rgb_resampler_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (pixel_rgb_resampler_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (pixel_rgb_resampler_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (pixel_rgb_resampler_avalon_rgb_source_data)           //                  .data
	);

	Video_System_Pixel_Scaler pixel_scaler (
		.clk                      (clock_signals_sys_clk_clk),                           //          clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                      //    clock_reset_reset.reset
		.stream_in_startofpacket  (pixel_rgb_resampler_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (pixel_rgb_resampler_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (pixel_rgb_resampler_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (pixel_rgb_resampler_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (pixel_rgb_resampler_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (pixel_scaler_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (pixel_scaler_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (pixel_scaler_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (pixel_scaler_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (pixel_scaler_avalon_scaler_source_data)               //                     .data
	);

	Video_System_VGA_Controller vga_controller (
		.clk           (clock_signals_vga_clk_clk),                             //        clock_reset.clk
		.reset         (rst_controller_001_reset_out_reset),                    //  clock_reset_reset.reset
		.data          (dual_clock_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (dual_clock_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (dual_clock_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (VGA_CLK_from_the_VGA_Controller),                       // external_interface.export
		.VGA_HS        (VGA_HS_from_the_VGA_Controller),                        //                   .export
		.VGA_VS        (VGA_VS_from_the_VGA_Controller),                        //                   .export
		.VGA_BLANK     (VGA_BLANK_from_the_VGA_Controller),                     //                   .export
		.VGA_SYNC      (VGA_SYNC_from_the_VGA_Controller),                      //                   .export
		.VGA_R         (VGA_R_from_the_VGA_Controller),                         //                   .export
		.VGA_G         (VGA_G_from_the_VGA_Controller),                         //                   .export
		.VGA_B         (VGA_B_from_the_VGA_Controller)                          //                   .export
	);

	Video_System_Video_In_Decoder video_in_decoder (
		.clk                      (clock_signals_sys_clk_clk),                            //           clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                       //     clock_reset_reset.reset
		.stream_out_ready         (video_in_decoder_avalon_decoder_source_ready),         // avalon_decoder_source.ready
		.stream_out_startofpacket (video_in_decoder_avalon_decoder_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (video_in_decoder_avalon_decoder_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (video_in_decoder_avalon_decoder_source_valid),         //                      .valid
		.stream_out_data          (video_in_decoder_avalon_decoder_source_data),          //                      .data
		.PIXEL_CLK                (Video_In_Decoder_external_interface_PIXEL_CLK),        //    external_interface.export
		.LINE_VALID               (Video_In_Decoder_external_interface_LINE_VALID),       //                      .export
		.FRAME_VALID              (Video_In_Decoder_external_interface_FRAME_VALID),      //                      .export
		.pixel_clk_reset          (Video_In_Decoder_external_interface_pixel_clk_reset),  //                      .export
		.PIXEL_DATA               (Video_In_Decoder_external_interface_PIXEL_DATA)        //                      .export
	);

	Video_System_Video_RGB_Resampler video_rgb_resampler (
		.clk                      (clock_signals_sys_clk_clk),                            //       clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                       // clock_reset_reset.reset
		.stream_in_startofpacket  (video_in_decoder_avalon_decoder_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (video_in_decoder_avalon_decoder_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (video_in_decoder_avalon_decoder_source_valid),         //                  .valid
		.stream_in_ready          (video_in_decoder_avalon_decoder_source_ready),         //                  .ready
		.stream_in_data           (video_in_decoder_avalon_decoder_source_data),          //                  .data
		.stream_out_ready         (video_rgb_resampler_avalon_rgb_source_ready),          // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_avalon_rgb_source_startofpacket),  //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_avalon_rgb_source_endofpacket),    //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_avalon_rgb_source_valid),          //                  .valid
		.stream_out_data          (video_rgb_resampler_avalon_rgb_source_data)            //                  .data
	);

	Video_System_Video_Clipper video_clipper (
		.clk                      (clock_signals_sys_clk_clk),                           //           clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                      //     clock_reset_reset.reset
		.stream_in_data           (video_rgb_resampler_avalon_rgb_source_data),          //   avalon_clipper_sink.data
		.stream_in_startofpacket  (video_rgb_resampler_avalon_rgb_source_startofpacket), //                      .startofpacket
		.stream_in_endofpacket    (video_rgb_resampler_avalon_rgb_source_endofpacket),   //                      .endofpacket
		.stream_in_valid          (video_rgb_resampler_avalon_rgb_source_valid),         //                      .valid
		.stream_in_ready          (video_rgb_resampler_avalon_rgb_source_ready),         //                      .ready
		.stream_out_ready         (video_clipper_avalon_clipper_source_ready),           // avalon_clipper_source.ready
		.stream_out_data          (video_clipper_avalon_clipper_source_data),            //                      .data
		.stream_out_startofpacket (video_clipper_avalon_clipper_source_startofpacket),   //                      .startofpacket
		.stream_out_endofpacket   (video_clipper_avalon_clipper_source_endofpacket),     //                      .endofpacket
		.stream_out_valid         (video_clipper_avalon_clipper_source_valid)            //                      .valid
	);

	Video_System_Video_Scaler video_scaler (
		.clk                      (clock_signals_sys_clk_clk),                         //          clock_reset.clk
		.reset                    (rst_controller_reset_out_reset),                    //    clock_reset_reset.reset
		.stream_in_startofpacket  (video_clipper_avalon_clipper_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (video_clipper_avalon_clipper_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (video_clipper_avalon_clipper_source_valid),         //                     .valid
		.stream_in_ready          (video_clipper_avalon_clipper_source_ready),         //                     .ready
		.stream_in_data           (video_clipper_avalon_clipper_source_data),          //                     .data
		.stream_out_ready         (video_scaler_avalon_scaler_source_ready),           // avalon_scaler_source.ready
		.stream_out_startofpacket (video_scaler_avalon_scaler_source_startofpacket),   //                     .startofpacket
		.stream_out_endofpacket   (video_scaler_avalon_scaler_source_endofpacket),     //                     .endofpacket
		.stream_out_valid         (video_scaler_avalon_scaler_source_valid),           //                     .valid
		.stream_out_data          (video_scaler_avalon_scaler_source_data)             //                     .data
	);

	Video_System_Video_DMA video_dma (
		.clk                  (clock_signals_sys_clk_clk),                                                    //              clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                                               //        clock_reset_reset.reset
		.stream_data          (video_scaler_avalon_scaler_source_data),                                       //          avalon_dma_sink.data
		.stream_startofpacket (video_scaler_avalon_scaler_source_startofpacket),                              //                         .startofpacket
		.stream_endofpacket   (video_scaler_avalon_scaler_source_endofpacket),                                //                         .endofpacket
		.stream_valid         (video_scaler_avalon_scaler_source_valid),                                      //                         .valid
		.stream_ready         (video_scaler_avalon_scaler_source_ready),                                      //                         .ready
		.slave_address        (video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable), //                         .byteenable
		.slave_read           (video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_read),       //                         .read
		.slave_write          (video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_write),      //                         .write
		.slave_writedata      (video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata),  //                         .writedata
		.slave_readdata       (video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata),   //                         .readdata
		.master_address       (video_dma_avalon_dma_master_address),                                          //        avalon_dma_master.address
		.master_waitrequest   (video_dma_avalon_dma_master_waitrequest),                                      //                         .waitrequest
		.master_write         (video_dma_avalon_dma_master_write),                                            //                         .write
		.master_writedata     (video_dma_avalon_dma_master_writedata)                                         //                         .writedata
	);

	Video_System_AV_Config av_config (
		.clk         (clock_signals_sys_clk_clk),                                                   //            clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                              //      clock_reset_reset.reset
		.address     (av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_address),     // avalon_av_config_slave.address
		.byteenable  (av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),  //                       .byteenable
		.read        (av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_read),        //                       .read
		.write       (av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_write),       //                       .write
		.writedata   (av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),   //                       .writedata
		.readdata    (av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),    //                       .readdata
		.waitrequest (av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest), //                       .waitrequest
		.I2C_SDAT    (I2C_SDAT_to_and_from_the_AV_Config),                                          //     external_interface.export
		.I2C_SCLK    (I2C_SCLK_from_the_AV_Config)                                                  //                       .export
	);

	Video_System_CPU cpu (
		.clk                                   (clock_signals_sys_clk_clk),                                          //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                    //                   reset_n.reset_n
		.d_address                             (cpu_data_master_address),                                            //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (cpu_data_master_read),                                               //                          .read
		.d_readdata                            (cpu_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (cpu_data_master_write),                                              //                          .write
		.d_writedata                           (cpu_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                                        //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                                 //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	Video_System_Clock_Signals clock_signals (
		.CLOCK_50    (clk),                                //       clk_in_primary.clk
		.reset       (rst_controller_002_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (clock_signals_sys_clk_clk),          //              sys_clk.clk
		.sys_reset_n (),                                   //        sys_clk_reset.reset_n
		.VGA_CLK     (clock_signals_vga_clk_clk)           //              vga_clk.clk
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (22),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_instruction_master_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                 //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address           (cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount         (1'b1),                                                                      //               (terminated)
		.av_byteenable         (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                      //               (terminated)
		.av_begintransfer      (1'b0),                                                                      //               (terminated)
		.av_chipselect         (1'b0),                                                                      //               (terminated)
		.av_readdatavalid      (),                                                                          //               (terminated)
		.av_write              (1'b0),                                                                      //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                      //               (terminated)
		.av_lock               (1'b0),                                                                      //               (terminated)
		.av_debugaccess        (1'b0),                                                                      //               (terminated)
		.uav_clken             (),                                                                          //               (terminated)
		.av_clken              (1'b1)                                                                       //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (22),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) cpu_data_master_translator (
		.clk                   (clock_signals_sys_clk_clk),                                          //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                     reset.reset
		.uav_address           (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_data_master_read),                                               //                          .read
		.av_readdata           (cpu_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_data_master_write),                                              //                          .write
		.av_writedata          (cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_readdatavalid      (),                                                                   //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) pixel_buffer_dma_avalon_pixel_dma_master_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                                   //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                              //                     reset.reset
		.uav_address           (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (pixel_buffer_dma_avalon_pixel_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),                                        //                          .waitrequest
		.av_read               (pixel_buffer_dma_avalon_pixel_dma_master_read),                                               //                          .read
		.av_readdata           (pixel_buffer_dma_avalon_pixel_dma_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),                                      //                          .readdatavalid
		.av_lock               (pixel_buffer_dma_avalon_pixel_dma_master_lock),                                               //                          .lock
		.av_burstcount         (1'b1),                                                                                        //               (terminated)
		.av_byteenable         (2'b11),                                                                                       //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                                        //               (terminated)
		.av_write              (1'b0),                                                                                        //               (terminated)
		.av_writedata          (16'b0000000000000000),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                                        //               (terminated)
		.uav_clken             (),                                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) video_dma_avalon_dma_master_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                      //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                     reset.reset
		.uav_address           (video_dma_avalon_dma_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (video_dma_avalon_dma_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (video_dma_avalon_dma_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (video_dma_avalon_dma_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (video_dma_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (video_dma_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (video_dma_avalon_dma_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (video_dma_avalon_dma_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (video_dma_avalon_dma_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (video_dma_avalon_dma_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (video_dma_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (video_dma_avalon_dma_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (video_dma_avalon_dma_master_waitrequest),                                        //                          .waitrequest
		.av_write              (video_dma_avalon_dma_master_write),                                              //                          .write
		.av_writedata          (video_dma_avalon_dma_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                           //               (terminated)
		.av_byteenable         (2'b11),                                                                          //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                           //               (terminated)
		.av_begintransfer      (1'b0),                                                                           //               (terminated)
		.av_chipselect         (1'b0),                                                                           //               (terminated)
		.av_read               (1'b0),                                                                           //               (terminated)
		.av_readdata           (),                                                                               //               (terminated)
		.av_readdatavalid      (),                                                                               //               (terminated)
		.av_lock               (1'b0),                                                                           //               (terminated)
		.av_debugaccess        (1'b0),                                                                           //               (terminated)
		.uav_clken             (),                                                                               //               (terminated)
		.av_clken              (1'b1)                                                                            //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_jtag_debug_module_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                   //                    reset.reset
		.uav_address           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (cpu_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                 //              (terminated)
		.av_lock               (),                                                                                 //              (terminated)
		.av_clken              (),                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                             //              (terminated)
		.av_outputenable       ()                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (12),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory_s1_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                   //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (onchip_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (onchip_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (onchip_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (onchip_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (onchip_memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (onchip_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (onchip_memory_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (20),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pixel_buffer_avalon_sram_slave_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (pixel_buffer_avalon_sram_slave_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_begintransfer      (),                                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                                          //              (terminated)
		.av_burstcount         (),                                                                                          //              (terminated)
		.av_waitrequest        (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                                          //              (terminated)
		.av_lock               (),                                                                                          //              (terminated)
		.av_chipselect         (),                                                                                          //              (terminated)
		.av_clken              (),                                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                                      //              (terminated)
		.av_debugaccess        (),                                                                                          //              (terminated)
		.av_outputenable       ()                                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) av_config_avalon_av_config_slave_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                              //                    reset.reset
		.uav_address           (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (av_config_avalon_av_config_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                                            //              (terminated)
		.av_burstcount         (),                                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                                            //              (terminated)
		.av_lock               (),                                                                                            //              (terminated)
		.av_chipselect         (),                                                                                            //              (terminated)
		.av_clken              (),                                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                                        //              (terminated)
		.av_debugaccess        (),                                                                                            //              (terminated)
		.av_outputenable       ()                                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) video_dma_avalon_dma_control_slave_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                //                    reset.reset
		.uav_address           (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (video_dma_avalon_dma_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer      (),                                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                                              //              (terminated)
		.av_burstcount         (),                                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                          //              (terminated)
		.av_waitrequest        (1'b0),                                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                                              //              (terminated)
		.av_lock               (),                                                                                              //              (terminated)
		.av_chipselect         (),                                                                                              //              (terminated)
		.av_clken              (),                                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                                          //              (terminated)
		.av_debugaccess        (),                                                                                              //              (terminated)
		.av_outputenable       ()                                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pixel_buffer_dma_avalon_control_slave_translator (
		.clk                   (clock_signals_sys_clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                   //                    reset.reset
		.uav_address           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (pixel_buffer_dma_avalon_control_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer      (),                                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                             //              (terminated)
		.av_waitrequest        (1'b0),                                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                                 //              (terminated)
		.av_lock               (),                                                                                                 //              (terminated)
		.av_chipselect         (),                                                                                                 //              (terminated)
		.av_clken              (),                                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                                  //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3)
	) cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clock_signals_sys_clk_clk),                                                          //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address       (cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                              //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                               //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                            //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                        //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                               //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clock_signals_sys_clk_clk),                                                   //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.av_address       (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                   //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                    //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                 //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                           //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                             //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                    //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.PKT_BEGIN_BURST           (61),
		.PKT_BURSTWRAP_H           (60),
		.PKT_BURSTWRAP_L           (58),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (55),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (64),
		.PKT_SRC_ID_L              (62),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (65),
		.ST_DATA_W                 (69),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (3),
		.BURSTWRAP_VALUE           (7)
	) pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent (
		.clk              (clock_signals_sys_clk_clk),                                                                            //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                                       // clk_reset.reset
		.av_address       (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_002_rsp_src_valid),                                                                            //        rp.valid
		.rp_data          (limiter_002_rsp_src_data),                                                                             //          .data
		.rp_channel       (limiter_002_rsp_src_channel),                                                                          //          .channel
		.rp_startofpacket (limiter_002_rsp_src_startofpacket),                                                                    //          .startofpacket
		.rp_endofpacket   (limiter_002_rsp_src_endofpacket),                                                                      //          .endofpacket
		.rp_ready         (limiter_002_rsp_src_ready)                                                                             //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.PKT_BEGIN_BURST           (61),
		.PKT_BURSTWRAP_H           (60),
		.PKT_BURSTWRAP_L           (58),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (55),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (64),
		.PKT_SRC_ID_L              (62),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (65),
		.ST_DATA_W                 (69),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (4),
		.BURSTWRAP_VALUE           (7)
	) video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent (
		.clk              (clock_signals_sys_clk_clk),                                                               //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.av_address       (video_dma_avalon_dma_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (video_dma_avalon_dma_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (video_dma_avalon_dma_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (video_dma_avalon_dma_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (video_dma_avalon_dma_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (video_dma_avalon_dma_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (video_dma_avalon_dma_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (video_dma_avalon_dma_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (video_dma_avalon_dma_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (video_dma_avalon_dma_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (video_dma_avalon_dma_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_003_rsp_src_valid),                                                               //        rp.valid
		.rp_data          (limiter_003_rsp_src_data),                                                                //          .data
		.rp_channel       (limiter_003_rsp_src_channel),                                                             //          .channel
		.rp_startofpacket (limiter_003_rsp_src_startofpacket),                                                       //          .startofpacket
		.rp_endofpacket   (limiter_003_rsp_src_endofpacket),                                                         //          .endofpacket
		.rp_ready         (limiter_003_rsp_src_ready)                                                                //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_signals_sys_clk_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                   //                .channel
		.rf_sink_ready           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_signals_sys_clk_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) onchip_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_signals_sys_clk_clk),                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                          //                .channel
		.rf_sink_ready           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_signals_sys_clk_clk),                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (61),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (64),
		.PKT_SRC_ID_L              (62),
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (65),
		.PKT_BURSTWRAP_H           (60),
		.PKT_BURSTWRAP_L           (58),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (55),
		.PKT_PROTECTION_H          (68),
		.PKT_PROTECTION_L          (68),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (69),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_signals_sys_clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                                         //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                                         //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                                          //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                                       //                .channel
		.rf_sink_ready           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (70),
		.FIFO_DEPTH          (3),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_signals_sys_clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_signals_sys_clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                        //       clk_reset.reset
		.m0_address              (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                                       //                .channel
		.rf_sink_ready           (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_signals_sys_clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                        // clk_reset.reset
		.in_data           (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                                  // (terminated)
		.csr_readdata      (),                                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                  // (terminated)
		.almost_full_data  (),                                                                                                      // (terminated)
		.almost_empty_data (),                                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                                  // (terminated)
		.out_empty         (),                                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                                  // (terminated)
		.out_error         (),                                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                                  // (terminated)
		.out_channel       ()                                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_signals_sys_clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                          //       clk_reset.reset
		.m0_address              (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                                         //                .channel
		.rf_sink_ready           (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_signals_sys_clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                          // clk_reset.reset
		.in_data           (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                                    // (terminated)
		.csr_readdata      (),                                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                    // (terminated)
		.almost_full_data  (),                                                                                                        // (terminated)
		.almost_empty_data (),                                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                                    // (terminated)
		.out_empty         (),                                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                                    // (terminated)
		.out_error         (),                                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                                    // (terminated)
		.out_channel       ()                                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_signals_sys_clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                             //       clk_reset.reset
		.m0_address              (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                                            //                .channel
		.rf_sink_ready           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_signals_sys_clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                             // clk_reset.reset
		.in_data           (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                                       // (terminated)
		.csr_readdata      (),                                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                       // (terminated)
		.almost_full_data  (),                                                                                                           // (terminated)
		.almost_empty_data (),                                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                                       // (terminated)
		.out_empty         (),                                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                                       // (terminated)
		.out_error         (),                                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                                       // (terminated)
		.out_channel       ()                                                                                                            // (terminated)
	);

	Video_System_addr_router addr_router (
		.sink_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                                              //          .valid
		.src_data           (addr_router_src_data),                                                               //          .data
		.src_channel        (addr_router_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                         //          .endofpacket
	);

	Video_System_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                   //          .valid
		.src_data           (addr_router_001_src_data),                                                    //          .data
		.src_channel        (addr_router_001_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                              //          .endofpacket
	);

	Video_System_addr_router_002 addr_router_002 (
		.sink_ready         (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pixel_buffer_dma_avalon_pixel_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                       // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                                            //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                                            //          .valid
		.src_data           (addr_router_002_src_data),                                                                             //          .data
		.src_channel        (addr_router_002_src_channel),                                                                          //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                                    //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                                       //          .endofpacket
	);

	Video_System_addr_router_002 addr_router_003 (
		.sink_ready         (video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (video_dma_avalon_dma_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                               //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                               //          .valid
		.src_data           (addr_router_003_src_data),                                                                //          .data
		.src_channel        (addr_router_003_src_channel),                                                             //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                          //          .endofpacket
	);

	Video_System_id_router id_router (
		.sink_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                              //       src.ready
		.src_valid          (id_router_src_valid),                                                              //          .valid
		.src_data           (id_router_src_data),                                                               //          .data
		.src_channel        (id_router_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                         //          .endofpacket
	);

	Video_System_id_router id_router_001 (
		.sink_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                     //       src.ready
		.src_valid          (id_router_001_src_valid),                                                     //          .valid
		.src_data           (id_router_001_src_data),                                                      //          .data
		.src_channel        (id_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                //          .endofpacket
	);

	Video_System_id_router_002 id_router_002 (
		.sink_ready         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pixel_buffer_avalon_sram_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                   //          .valid
		.src_data           (id_router_002_src_data),                                                                    //          .data
		.src_channel        (id_router_002_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                              //          .endofpacket
	);

	Video_System_id_router_003 id_router_003 (
		.sink_ready         (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (av_config_avalon_av_config_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                     //          .valid
		.src_data           (id_router_003_src_data),                                                                      //          .data
		.src_channel        (id_router_003_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                                //          .endofpacket
	);

	Video_System_id_router_003 id_router_004 (
		.sink_ready         (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (video_dma_avalon_dma_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                                       //       src.ready
		.src_valid          (id_router_004_src_valid),                                                                       //          .valid
		.src_data           (id_router_004_src_data),                                                                        //          .data
		.src_channel        (id_router_004_src_channel),                                                                     //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                                  //          .endofpacket
	);

	Video_System_id_router_003 id_router_005 (
		.sink_ready         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pixel_buffer_dma_avalon_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_signals_sys_clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                          //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                          //          .valid
		.src_data           (id_router_005_src_data),                                                                           //          .data
		.src_channel        (id_router_005_src_channel),                                                                        //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                                     //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (5),
		.PIPELINED                 (0),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (6),
		.VALID_WIDTH               (6),
		.ENFORCE_ORDER             (0),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clock_signals_sys_clk_clk),      //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (8),
		.PIPELINED                 (0),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (6),
		.VALID_WIDTH               (6),
		.ENFORCE_ORDER             (0),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clock_signals_sys_clk_clk),          //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (65),
		.PKT_TRANS_POSTED          (51),
		.MAX_OUTSTANDING_RESPONSES (8),
		.PIPELINED                 (0),
		.ST_DATA_W                 (69),
		.ST_CHANNEL_W              (6),
		.VALID_WIDTH               (6),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (55),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16)
	) limiter_002 (
		.clk                    (clock_signals_sys_clk_clk),             //       clk.clk
		.reset                  (rst_controller_reset_out_reset),        // clk_reset.reset
		.cmd_sink_ready         (addr_router_002_src_ready),             //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_002_src_valid),             //          .valid
		.cmd_sink_data          (addr_router_002_src_data),              //          .data
		.cmd_sink_channel       (addr_router_002_src_channel),           //          .channel
		.cmd_sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.cmd_src_ready          (limiter_002_cmd_src_ready),             //   cmd_src.ready
		.cmd_src_data           (limiter_002_cmd_src_data),              //          .data
		.cmd_src_channel        (limiter_002_cmd_src_channel),           //          .channel
		.cmd_src_startofpacket  (limiter_002_cmd_src_startofpacket),     //          .startofpacket
		.cmd_src_endofpacket    (limiter_002_cmd_src_endofpacket),       //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_demux_002_src1_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_002_rsp_src_ready),             //   rsp_src.ready
		.rsp_src_valid          (limiter_002_rsp_src_valid),             //          .valid
		.rsp_src_data           (limiter_002_rsp_src_data),              //          .data
		.rsp_src_channel        (limiter_002_rsp_src_channel),           //          .channel
		.rsp_src_startofpacket  (limiter_002_rsp_src_startofpacket),     //          .startofpacket
		.rsp_src_endofpacket    (limiter_002_rsp_src_endofpacket),       //          .endofpacket
		.cmd_src_valid          (limiter_002_cmd_valid_data)             // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (67),
		.PKT_DEST_ID_L             (65),
		.PKT_TRANS_POSTED          (51),
		.MAX_OUTSTANDING_RESPONSES (8),
		.PIPELINED                 (0),
		.ST_DATA_W                 (69),
		.ST_CHANNEL_W              (6),
		.VALID_WIDTH               (6),
		.ENFORCE_ORDER             (0),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (55),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16)
	) limiter_003 (
		.clk                    (clock_signals_sys_clk_clk),             //       clk.clk
		.reset                  (rst_controller_reset_out_reset),        // clk_reset.reset
		.cmd_sink_ready         (addr_router_003_src_ready),             //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_003_src_valid),             //          .valid
		.cmd_sink_data          (addr_router_003_src_data),              //          .data
		.cmd_sink_channel       (addr_router_003_src_channel),           //          .channel
		.cmd_sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.cmd_src_ready          (limiter_003_cmd_src_ready),             //   cmd_src.ready
		.cmd_src_data           (limiter_003_cmd_src_data),              //          .data
		.cmd_src_channel        (limiter_003_cmd_src_channel),           //          .channel
		.cmd_src_startofpacket  (limiter_003_cmd_src_startofpacket),     //          .startofpacket
		.cmd_src_endofpacket    (limiter_003_cmd_src_endofpacket),       //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_demux_002_src2_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_demux_002_src2_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_demux_002_src2_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_demux_002_src2_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_003_rsp_src_ready),             //   rsp_src.ready
		.rsp_src_valid          (limiter_003_rsp_src_valid),             //          .valid
		.rsp_src_data           (limiter_003_rsp_src_data),              //          .data
		.rsp_src_channel        (limiter_003_rsp_src_channel),           //          .channel
		.rsp_src_startofpacket  (limiter_003_rsp_src_startofpacket),     //          .startofpacket
		.rsp_src_endofpacket    (limiter_003_rsp_src_endofpacket),       //          .endofpacket
		.cmd_src_valid          (limiter_003_cmd_valid_data)             // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (61),
		.PKT_BYTE_CNT_H            (57),
		.PKT_BYTE_CNT_L            (55),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURSTWRAP_H           (60),
		.PKT_BURSTWRAP_L           (58),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.ST_DATA_W                 (69),
		.ST_CHANNEL_W              (6),
		.OUT_BYTE_CNT_H            (56),
		.OUT_BURSTWRAP_H           (60),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter (
		.clk                   (clock_signals_sys_clk_clk),           //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_002_src_valid),          //     sink0.valid
		.sink0_data            (cmd_xbar_mux_002_src_data),           //          .data
		.sink0_channel         (cmd_xbar_mux_002_src_channel),        //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_002_src_startofpacket),  //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_002_src_endofpacket),    //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_002_src_ready),          //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_n),                          // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clock_signals_sys_clk_clk),         //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_in2  (1'b0),                              // (terminated)
		.reset_in3  (1'b0),                              // (terminated)
		.reset_in4  (1'b0),                              // (terminated)
		.reset_in5  (1'b0),                              // (terminated)
		.reset_in6  (1'b0),                              // (terminated)
		.reset_in7  (1'b0),                              // (terminated)
		.reset_in8  (1'b0),                              // (terminated)
		.reset_in9  (1'b0),                              // (terminated)
		.reset_in10 (1'b0),                              // (terminated)
		.reset_in11 (1'b0),                              // (terminated)
		.reset_in12 (1'b0),                              // (terminated)
		.reset_in13 (1'b0),                              // (terminated)
		.reset_in14 (1'b0),                              // (terminated)
		.reset_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk        (clock_signals_vga_clk_clk),          //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (cpu_jtag_debug_module_reset_reset),  // reset_in0.reset
		.reset_in1  (~reset_n),                           // reset_in1.reset
		.clk        (clk),                                //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	Video_System_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clock_signals_sys_clk_clk),         //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //           .endofpacket
	);

	Video_System_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clock_signals_sys_clk_clk),             //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket)    //           .endofpacket
	);

	Video_System_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (clock_signals_sys_clk_clk),             //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_002_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_002_cmd_src_channel),           //           .channel
		.sink_data          (limiter_002_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_002_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_002_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_002_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //           .endofpacket
	);

	Video_System_cmd_xbar_demux_002 cmd_xbar_demux_003 (
		.clk                (clock_signals_sys_clk_clk),             //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_003_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_003_cmd_src_channel),           //           .channel
		.sink_data          (limiter_003_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_003_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_003_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_003_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //           .endofpacket
	);

	Video_System_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clock_signals_sys_clk_clk),             //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	Video_System_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clock_signals_sys_clk_clk),             //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	Video_System_cmd_xbar_mux_002 cmd_xbar_mux_002 (
		.clk                 (clock_signals_sys_clk_clk),             //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_src_ready),               //     sink0.ready
		.sink0_valid         (width_adapter_src_valid),               //          .valid
		.sink0_channel       (width_adapter_src_channel),             //          .channel
		.sink0_data          (width_adapter_src_data),                //          .data
		.sink0_startofpacket (width_adapter_src_startofpacket),       //          .startofpacket
		.sink0_endofpacket   (width_adapter_src_endofpacket),         //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_003_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	Video_System_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clock_signals_sys_clk_clk),         //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	Video_System_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clock_signals_sys_clk_clk),             //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	Video_System_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clock_signals_sys_clk_clk),             //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_002_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_002_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_002_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_002_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_002_src2_endofpacket)    //          .endofpacket
	);

	Video_System_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (clock_signals_sys_clk_clk),             //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	Video_System_rsp_xbar_demux_003 rsp_xbar_demux_004 (
		.clk                (clock_signals_sys_clk_clk),             //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	Video_System_rsp_xbar_demux_003 rsp_xbar_demux_005 (
		.clk                (clock_signals_sys_clk_clk),             //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	Video_System_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clock_signals_sys_clk_clk),             //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	Video_System_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (clock_signals_sys_clk_clk),             //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (width_adapter_001_src_ready),           //     sink2.ready
		.sink2_valid         (width_adapter_001_src_valid),           //          .valid
		.sink2_channel       (width_adapter_001_src_channel),         //          .channel
		.sink2_data          (width_adapter_001_src_data),            //          .data
		.sink2_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink2_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (87),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (57),
		.OUT_PKT_BYTE_CNT_L            (55),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_ST_DATA_W                 (69),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk               (clock_signals_sys_clk_clk),             //       clk.clk
		.reset             (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid          (cmd_xbar_demux_001_src2_valid),         //      sink.valid
		.in_channel        (cmd_xbar_demux_001_src2_channel),       //          .channel
		.in_startofpacket  (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.in_ready          (cmd_xbar_demux_001_src2_ready),         //          .ready
		.in_data           (cmd_xbar_demux_001_src2_data),          //          .data
		.out_endofpacket   (width_adapter_src_endofpacket),         //       src.endofpacket
		.out_data          (width_adapter_src_data),                //          .data
		.out_channel       (width_adapter_src_channel),             //          .channel
		.out_valid         (width_adapter_src_valid),               //          .valid
		.out_ready         (width_adapter_src_ready),               //          .ready
		.out_startofpacket (width_adapter_src_startofpacket)        //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (57),
		.IN_PKT_BYTE_CNT_L             (55),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (60),
		.IN_PKT_BURSTWRAP_L            (58),
		.IN_ST_DATA_W                  (69),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (87),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk               (clock_signals_sys_clk_clk),             //       clk.clk
		.reset             (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid          (rsp_xbar_demux_002_src0_valid),         //      sink.valid
		.in_channel        (rsp_xbar_demux_002_src0_channel),       //          .channel
		.in_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.in_ready          (rsp_xbar_demux_002_src0_ready),         //          .ready
		.in_data           (rsp_xbar_demux_002_src0_data),          //          .data
		.out_endofpacket   (width_adapter_001_src_endofpacket),     //       src.endofpacket
		.out_data          (width_adapter_001_src_data),            //          .data
		.out_channel       (width_adapter_001_src_channel),         //          .channel
		.out_valid         (width_adapter_001_src_valid),           //          .valid
		.out_ready         (width_adapter_001_src_ready),           //          .ready
		.out_startofpacket (width_adapter_001_src_startofpacket)    //          .startofpacket
	);

	Video_System_irq_mapper irq_mapper (
		.clk        (clock_signals_sys_clk_clk),      //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (cpu_d_irq_irq)                   //    sender.irq
	);

endmodule
