module ZEXT(
	input logic [15:0] in,

	output logic [19:0] out
);

	assign out = in;

endmodule



